`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2016/01/29 23:04:25
// Design Name: 
// Module Name: notgate_sim
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module notgate_sim(

    );
    // input 
reg [31:0] a=32'h00000000;

//outbut
wire [31:0] c;
 notgate #(32) u(a,c);    // ʵ�������ŵ�ʱ���趨���Ϊ32

initial begin
#100  a=32'hffffffff;
#100  a=32'hf070ff5f;
end
endmodule
