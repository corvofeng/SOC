`timescale 1ns / 1ps
/*
 *=============================================================================
 *    Filename:input1.v
 *
 *     Version: 1.0
 *  Created on: July 11, 2016
 *    
 *      Author: corvo
 *=============================================================================
 */
 
module input0(
    zero
    );
    output[31:0] zero;
    assign zero = 32'h0;
endmodule
