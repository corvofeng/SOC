/*
 *=============================================================================
 *    Filename: alu_test.v
 *
 *     Version: 1.0
 *  Created on: September 19, 2017
 *
 *      Author: corvo
 *=============================================================================
 */


module alu_test();


    initial begin
        $display("Hello, World!");
        $finish;
    end

endmodule

