`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2017/09/25 14:54:17
// Design Name:
// Module Name: pc_sim
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module pc_sim(

       );
//    reg clk,clrn;
//    wire [31:0]ins,bpc,dpc,jpc,pc4,npc;
//    reg []
//    reg [1:0]pcsource;

//    socpc ipc(
//      .pc(pc),
//      .bpc(bpc),
//      .dpc(dpc),
//      .jpc(jpc),
//      .pcsource(pcsource),
//      .pc4(pc4),
//      .ins(ins),
//      .npc(npc)
//        );
//    initial begin
//          #1 clrn=1;
//             clk=0;
//             pcsource= 2'b00;
//          #5 clrn = 0;
//         #500 clrn = 1;
//           end
//           always #5 clk=~clk;

endmodule
